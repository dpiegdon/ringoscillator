
module top(input CLK, output J1_10);

	ringoscillator r0 (CLK, J1_10);

endmodule
