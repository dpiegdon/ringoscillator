
module top(input CLK, output J1_10);

	wire random;

	wire s0, s1, s2, s3;

	ringoscillator r0(s0);
	ringoscillator r1(s1);
	ringoscillator r2(s2);
	ringoscillator r3(s3);

	SB_LUT4 #(
		.LUT_INIT(16'b1010_1100_1110_0001)
	) buffers (
		.O(random),
		.I0(s0),
		.I1(s1),
		.I2(s2),
		.I3(s3)
	);

	wire [0:15] lfsr;
	lfsr_fibonacci fibo(CLK, 0, random, lfsr);

	assign J1_10 = lfsr[15];

endmodule
